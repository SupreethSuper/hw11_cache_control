localparam ALU_PASS1 = 4'h0;
localparam ALU_ADD   = 4'h1;
localparam ALU_AND   = 4'h2;
localparam ALU_OR    = 4'h3;
localparam ALU_NOR   = 4'h4;
localparam ALU_SUB   = 4'h5;
localparam ALU_LTS   = 4'h6;
localparam ALU_LTU   = 4'h7;
localparam ALU_SLL   = 4'h8;
localparam ALU_SRL   = 4'h9;
localparam ALU_PASS2 = 4'hA;
localparam ALU_SRA   = 4'hB;
